NOR2 Simulation
.lib "/usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt

.param theWidth = 650000u

* NOR2 Gate
X0 NODO A VPWR NWELL sky130_fd_pr__pfet_01v8 w={theWidth} l=150000u
X1 Y    B NODO NWELL sky130_fd_pr__pfet_01v8 w={theWidth} l=150000u

X2 Y A VGND VSUBS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND B Y VSUBS sky130_fd_pr__nfet_01v8 w=650000u l=150000u

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create pulse
Va A VGND pulse(0 1.8 1p 10p 10p 2n 4n)
Vb B VGND pulse(0 1.8 1p 10p 10p 1n 2n)
.tran 10e-12 4e-09 0e-00

.control 
    let runs = 20
    let i = 0
    set c = " "
    dowhile i < runs
      let newp = 600000u + i * 50000u
      alterparam theWidth = $&newp
      reset
      run
      let i = i + 1
    end
    let j = 1
    dowhile j <= runs
      set c = ( $c tran{$&j}.Y )
      let j = j + 1
    end
    plot A+4 B+2 $c xlabel "Time [ns]" ylabel "Voltage [V]"  title "NOR2 Gate optimization"
    plot tran1.Y tran10.Y tran5.Y
*   quit
.endc

.end
