NOR2 Simulation
.lib "/usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt


X0 NODO A VPWR VPWR sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X1 Y    B NODO VPWR sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u

X2 Y A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND B Y VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u


* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create pulse
Va A VGND pulse(0 1.8 1p 10p 10p 2n 4n)
Vb B VGND pulse(0 1.8 1p 10p 10p 1n 2n)
.tran 10e-12 4e-09 0e-00

.control
run
set color0 = white
set color1 = black
plot A+2 B Y-2
plot i(Vdd)
.endc

.end
